// PCIe_rsa.v

// Generated using ACDS version 14.1 186 at 2015.05.05.20:21:05

`timescale 1 ps / 1 ps
module PCIe_rsa (
		input  wire [31:0] avalon_shell_rsa_0_m0_address_address,         //     avalon_shell_rsa_0_m0_address.address
		input  wire        avalon_shell_rsa_0_m0_read_read,               //        avalon_shell_rsa_0_m0_read.read
		output wire [7:0]  avalon_shell_rsa_0_m0_readdata_readdata,       //    avalon_shell_rsa_0_m0_readdata.readdata
		output wire        avalon_shell_rsa_0_m0_waitrequest_waitrequest, // avalon_shell_rsa_0_m0_waitrequest.waitrequest
		input  wire        avalon_shell_rsa_0_m0_write_write,             //       avalon_shell_rsa_0_m0_write.write
		input  wire [7:0]  avalon_shell_rsa_0_m0_writedata_writedata,     //   avalon_shell_rsa_0_m0_writedata.writedata
		output wire        avalon_shell_rsa_0_s0_address_address,         //     avalon_shell_rsa_0_s0_address.address
		output wire        avalon_shell_rsa_0_s0_read_read,               //        avalon_shell_rsa_0_s0_read.read
		input  wire [7:0]  avalon_shell_rsa_0_s0_readdata_readdata,       //    avalon_shell_rsa_0_s0_readdata.readdata
		input  wire        avalon_shell_rsa_0_s0_waitrequest_waitrequest, // avalon_shell_rsa_0_s0_waitrequest.waitrequest
		output wire        avalon_shell_rsa_0_s0_write_write,             //       avalon_shell_rsa_0_s0_write.write
		output wire [7:0]  avalon_shell_rsa_0_s0_writedata_writedata,     //   avalon_shell_rsa_0_s0_writedata.writedata
		input  wire        clk_0_clk,                                     //                             clk_0.clk
		output wire [14:0] ddr3a_mem_a,                                   //                             ddr3a.mem_a
		output wire [2:0]  ddr3a_mem_ba,                                  //                                  .mem_ba
		output wire [0:0]  ddr3a_mem_ck,                                  //                                  .mem_ck
		output wire [0:0]  ddr3a_mem_ck_n,                                //                                  .mem_ck_n
		output wire [0:0]  ddr3a_mem_cke,                                 //                                  .mem_cke
		output wire [0:0]  ddr3a_mem_cs_n,                                //                                  .mem_cs_n
		output wire [7:0]  ddr3a_mem_dm,                                  //                                  .mem_dm
		output wire [0:0]  ddr3a_mem_ras_n,                               //                                  .mem_ras_n
		output wire [0:0]  ddr3a_mem_cas_n,                               //                                  .mem_cas_n
		output wire [0:0]  ddr3a_mem_we_n,                                //                                  .mem_we_n
		output wire        ddr3a_mem_reset_n,                             //                                  .mem_reset_n
		inout  wire [63:0] ddr3a_mem_dq,                                  //                                  .mem_dq
		inout  wire [7:0]  ddr3a_mem_dqs,                                 //                                  .mem_dqs
		inout  wire [7:0]  ddr3a_mem_dqs_n,                               //                                  .mem_dqs_n
		output wire [0:0]  ddr3a_mem_odt,                                 //                                  .mem_odt
		input  wire        ddr3a_oct_rzqin,                               //                         ddr3a_oct.rzqin
		output wire        ddr3a_pll_sharing_pll_mem_clk,                 //                 ddr3a_pll_sharing.pll_mem_clk
		output wire        ddr3a_pll_sharing_pll_write_clk,               //                                  .pll_write_clk
		output wire        ddr3a_pll_sharing_pll_locked,                  //                                  .pll_locked
		output wire        ddr3a_pll_sharing_pll_write_clk_pre_phy_clk,   //                                  .pll_write_clk_pre_phy_clk
		output wire        ddr3a_pll_sharing_pll_addr_cmd_clk,            //                                  .pll_addr_cmd_clk
		output wire        ddr3a_pll_sharing_pll_avl_clk,                 //                                  .pll_avl_clk
		output wire        ddr3a_pll_sharing_pll_config_clk,              //                                  .pll_config_clk
		output wire        ddr3a_pll_sharing_pll_hr_clk,                  //                                  .pll_hr_clk
		output wire        ddr3a_pll_sharing_pll_p2c_read_clk,            //                                  .pll_p2c_read_clk
		output wire        ddr3a_pll_sharing_pll_c2p_write_clk,           //                                  .pll_c2p_write_clk
		output wire        ddr3a_status_local_init_done,                  //                      ddr3a_status.local_init_done
		output wire        ddr3a_status_local_cal_success,                //                                  .local_cal_success
		output wire        ddr3a_status_local_cal_fail,                   //                                  .local_cal_fail
		input  wire        pcie_interface_hip_serial_rx_in0,              //         pcie_interface_hip_serial.rx_in0
		input  wire        pcie_interface_hip_serial_rx_in1,              //                                  .rx_in1
		input  wire        pcie_interface_hip_serial_rx_in2,              //                                  .rx_in2
		input  wire        pcie_interface_hip_serial_rx_in3,              //                                  .rx_in3
		input  wire        pcie_interface_hip_serial_rx_in4,              //                                  .rx_in4
		input  wire        pcie_interface_hip_serial_rx_in5,              //                                  .rx_in5
		input  wire        pcie_interface_hip_serial_rx_in6,              //                                  .rx_in6
		input  wire        pcie_interface_hip_serial_rx_in7,              //                                  .rx_in7
		output wire        pcie_interface_hip_serial_tx_out0,             //                                  .tx_out0
		output wire        pcie_interface_hip_serial_tx_out1,             //                                  .tx_out1
		output wire        pcie_interface_hip_serial_tx_out2,             //                                  .tx_out2
		output wire        pcie_interface_hip_serial_tx_out3,             //                                  .tx_out3
		output wire        pcie_interface_hip_serial_tx_out4,             //                                  .tx_out4
		output wire        pcie_interface_hip_serial_tx_out5,             //                                  .tx_out5
		output wire        pcie_interface_hip_serial_tx_out6,             //                                  .tx_out6
		output wire        pcie_interface_hip_serial_tx_out7,             //                                  .tx_out7
		input  wire        pcie_interface_npor_npor,                      //               pcie_interface_npor.npor
		input  wire        pcie_interface_npor_pin_perst,                 //                                  .pin_perst
		input  wire        pcie_interface_refclk_clk,                     //             pcie_interface_refclk.clk
		input  wire        reset_0_reset_n                                //                           reset_0.reset_n
	);

	wire   [31:0] pcie_config_driver_reconfig_mgmt_readdata;            // PCIe_config:reconfig_mgmt_readdata -> PCIe_config_driver:reconfig_mgmt_readdata
	wire          pcie_config_driver_reconfig_mgmt_waitrequest;         // PCIe_config:reconfig_mgmt_waitrequest -> PCIe_config_driver:reconfig_mgmt_waitrequest
	wire    [6:0] pcie_config_driver_reconfig_mgmt_address;             // PCIe_config_driver:reconfig_mgmt_address -> PCIe_config:reconfig_mgmt_address
	wire          pcie_config_driver_reconfig_mgmt_read;                // PCIe_config_driver:reconfig_mgmt_read -> PCIe_config:reconfig_mgmt_read
	wire          pcie_config_driver_reconfig_mgmt_write;               // PCIe_config_driver:reconfig_mgmt_write -> PCIe_config:reconfig_mgmt_write
	wire   [31:0] pcie_config_driver_reconfig_mgmt_writedata;           // PCIe_config_driver:reconfig_mgmt_writedata -> PCIe_config:reconfig_mgmt_writedata
	wire          pcie_interface_coreclkout_clk;                        // PCIE_interface:coreclkout -> [PCIe_config_driver:pld_clk, dma0:clk, dma0_pp:clk, irq_mapper:clk, mm_interconnect_0:PCIE_interface_coreclkout_clk, mm_interconnect_1:PCIE_interface_coreclkout_clk, mm_interconnect_2:PCIE_interface_coreclkout_clk, mm_interconnect_3:PCIE_interface_coreclkout_clk, rst_controller_001:clk]
	wire    [1:0] pcie_interface_hip_currentspeed_currentspeed;         // PCIE_interface:currentspeed -> PCIe_config_driver:currentspeed
	wire          pcie_interface_hip_status_derr_cor_ext_rcv;           // PCIE_interface:derr_cor_ext_rcv -> PCIe_config_driver:derr_cor_ext_rcv_drv
	wire          pcie_interface_hip_status_hotrst_exit;                // PCIE_interface:hotrst_exit -> PCIe_config_driver:hotrst_exit_drv
	wire          pcie_interface_hip_status_rx_par_err;                 // PCIE_interface:rx_par_err -> PCIe_config_driver:rx_par_err_drv
	wire   [11:0] pcie_interface_hip_status_ko_cpl_spc_data;            // PCIE_interface:ko_cpl_spc_data -> PCIe_config_driver:ko_cpl_spc_data_drv
	wire          pcie_interface_hip_status_dlup_exit;                  // PCIE_interface:dlup_exit -> PCIe_config_driver:dlup_exit_drv
	wire          pcie_interface_hip_status_derr_cor_ext_rpl;           // PCIE_interface:derr_cor_ext_rpl -> PCIe_config_driver:derr_cor_ext_rpl_drv
	wire          pcie_interface_hip_status_l2_exit;                    // PCIE_interface:l2_exit -> PCIe_config_driver:l2_exit_drv
	wire          pcie_interface_hip_status_dlup;                       // PCIE_interface:dlup -> PCIe_config_driver:dlup_drv
	wire    [3:0] pcie_interface_hip_status_int_status;                 // PCIE_interface:int_status -> PCIe_config_driver:int_status_drv
	wire          pcie_interface_hip_status_ev128ns;                    // PCIE_interface:ev128ns -> PCIe_config_driver:ev128ns_drv
	wire    [4:0] pcie_interface_hip_status_ltssmstate;                 // PCIE_interface:ltssmstate -> PCIe_config_driver:ltssmstate_drv
	wire    [1:0] pcie_interface_hip_status_tx_par_err;                 // PCIE_interface:tx_par_err -> PCIe_config_driver:tx_par_err_drv
	wire    [3:0] pcie_interface_hip_status_lane_act;                   // PCIE_interface:lane_act -> PCIe_config_driver:lane_act_drv
	wire          pcie_interface_hip_status_cfg_par_err;                // PCIE_interface:cfg_par_err -> PCIe_config_driver:cfg_par_err_drv
	wire          pcie_interface_hip_status_derr_rpl;                   // PCIE_interface:derr_rpl -> PCIe_config_driver:derr_rpl_drv
	wire          pcie_interface_hip_status_ev1us;                      // PCIE_interface:ev1us -> PCIe_config_driver:ev1us_drv
	wire    [7:0] pcie_interface_hip_status_ko_cpl_spc_header;          // PCIE_interface:ko_cpl_spc_header -> PCIe_config_driver:ko_cpl_spc_header_drv
	wire          pcie_config_reconfig_busy_reconfig_busy;              // PCIe_config:reconfig_busy -> PCIe_config_driver:reconfig_busy
	wire  [459:0] pcie_interface_reconfig_from_xcvr_reconfig_from_xcvr; // PCIE_interface:reconfig_from_xcvr -> PCIe_config:reconfig_from_xcvr
	wire  [699:0] pcie_config_reconfig_to_xcvr_reconfig_to_xcvr;        // PCIe_config:reconfig_to_xcvr -> PCIE_interface:reconfig_to_xcvr
	wire          pcie_interface_rxm_bar0_waitrequest;                  // mm_interconnect_0:PCIE_interface_Rxm_BAR0_waitrequest -> PCIE_interface:RxmWaitRequest_0_i
	wire  [127:0] pcie_interface_rxm_bar0_readdata;                     // mm_interconnect_0:PCIE_interface_Rxm_BAR0_readdata -> PCIE_interface:RxmReadData_0_i
	wire   [31:0] pcie_interface_rxm_bar0_address;                      // PCIE_interface:RxmAddress_0_o -> mm_interconnect_0:PCIE_interface_Rxm_BAR0_address
	wire          pcie_interface_rxm_bar0_read;                         // PCIE_interface:RxmRead_0_o -> mm_interconnect_0:PCIE_interface_Rxm_BAR0_read
	wire   [15:0] pcie_interface_rxm_bar0_byteenable;                   // PCIE_interface:RxmByteEnable_0_o -> mm_interconnect_0:PCIE_interface_Rxm_BAR0_byteenable
	wire          pcie_interface_rxm_bar0_readdatavalid;                // mm_interconnect_0:PCIE_interface_Rxm_BAR0_readdatavalid -> PCIE_interface:RxmReadDataValid_0_i
	wire          pcie_interface_rxm_bar0_write;                        // PCIE_interface:RxmWrite_0_o -> mm_interconnect_0:PCIE_interface_Rxm_BAR0_write
	wire  [127:0] pcie_interface_rxm_bar0_writedata;                    // PCIE_interface:RxmWriteData_0_o -> mm_interconnect_0:PCIE_interface_Rxm_BAR0_writedata
	wire    [5:0] pcie_interface_rxm_bar0_burstcount;                   // PCIE_interface:RxmBurstCount_0_o -> mm_interconnect_0:PCIE_interface_Rxm_BAR0_burstcount
	wire          mm_interconnect_0_pcie_interface_cra_chipselect;      // mm_interconnect_0:PCIE_interface_Cra_chipselect -> PCIE_interface:CraChipSelect_i
	wire   [31:0] mm_interconnect_0_pcie_interface_cra_readdata;        // PCIE_interface:CraReadData_o -> mm_interconnect_0:PCIE_interface_Cra_readdata
	wire          mm_interconnect_0_pcie_interface_cra_waitrequest;     // PCIE_interface:CraWaitRequest_o -> mm_interconnect_0:PCIE_interface_Cra_waitrequest
	wire   [13:0] mm_interconnect_0_pcie_interface_cra_address;         // mm_interconnect_0:PCIE_interface_Cra_address -> PCIE_interface:CraAddress_i
	wire          mm_interconnect_0_pcie_interface_cra_read;            // mm_interconnect_0:PCIE_interface_Cra_read -> PCIE_interface:CraRead
	wire    [3:0] mm_interconnect_0_pcie_interface_cra_byteenable;      // mm_interconnect_0:PCIE_interface_Cra_byteenable -> PCIE_interface:CraByteEnable_i
	wire          mm_interconnect_0_pcie_interface_cra_write;           // mm_interconnect_0:PCIE_interface_Cra_write -> PCIE_interface:CraWrite
	wire   [31:0] mm_interconnect_0_pcie_interface_cra_writedata;       // mm_interconnect_0:PCIE_interface_Cra_writedata -> PCIE_interface:CraWriteData_i
	wire          mm_interconnect_0_dma0_control_port_slave_chipselect; // mm_interconnect_0:dma0_control_port_slave_chipselect -> dma0:dma_ctl_chipselect
	wire   [31:0] mm_interconnect_0_dma0_control_port_slave_readdata;   // dma0:dma_ctl_readdata -> mm_interconnect_0:dma0_control_port_slave_readdata
	wire    [2:0] mm_interconnect_0_dma0_control_port_slave_address;    // mm_interconnect_0:dma0_control_port_slave_address -> dma0:dma_ctl_address
	wire          mm_interconnect_0_dma0_control_port_slave_write;      // mm_interconnect_0:dma0_control_port_slave_write -> dma0:dma_ctl_write_n
	wire   [31:0] mm_interconnect_0_dma0_control_port_slave_writedata;  // mm_interconnect_0:dma0_control_port_slave_writedata -> dma0:dma_ctl_writedata
	wire          pcie_interface_rxm_bar2_waitrequest;                  // mm_interconnect_1:PCIE_interface_Rxm_BAR2_waitrequest -> PCIE_interface:RxmWaitRequest_2_i
	wire  [127:0] pcie_interface_rxm_bar2_readdata;                     // mm_interconnect_1:PCIE_interface_Rxm_BAR2_readdata -> PCIE_interface:RxmReadData_2_i
	wire   [31:0] pcie_interface_rxm_bar2_address;                      // PCIE_interface:RxmAddress_2_o -> mm_interconnect_1:PCIE_interface_Rxm_BAR2_address
	wire          pcie_interface_rxm_bar2_read;                         // PCIE_interface:RxmRead_2_o -> mm_interconnect_1:PCIE_interface_Rxm_BAR2_read
	wire   [15:0] pcie_interface_rxm_bar2_byteenable;                   // PCIE_interface:RxmByteEnable_2_o -> mm_interconnect_1:PCIE_interface_Rxm_BAR2_byteenable
	wire          pcie_interface_rxm_bar2_readdatavalid;                // mm_interconnect_1:PCIE_interface_Rxm_BAR2_readdatavalid -> PCIE_interface:RxmReadDataValid_2_i
	wire          pcie_interface_rxm_bar2_write;                        // PCIE_interface:RxmWrite_2_o -> mm_interconnect_1:PCIE_interface_Rxm_BAR2_write
	wire  [127:0] pcie_interface_rxm_bar2_writedata;                    // PCIE_interface:RxmWriteData_2_o -> mm_interconnect_1:PCIE_interface_Rxm_BAR2_writedata
	wire    [5:0] pcie_interface_rxm_bar2_burstcount;                   // PCIE_interface:RxmBurstCount_2_o -> mm_interconnect_1:PCIE_interface_Rxm_BAR2_burstcount
	wire  [127:0] mm_interconnect_1_avalon_shell_rsa_0_s0_readdata;     // avalon_shell_rsa_0:avs_s0_readdata -> mm_interconnect_1:avalon_shell_rsa_0_s0_readdata
	wire          mm_interconnect_1_avalon_shell_rsa_0_s0_waitrequest;  // avalon_shell_rsa_0:avs_s0_waitrequest -> mm_interconnect_1:avalon_shell_rsa_0_s0_waitrequest
	wire    [0:0] mm_interconnect_1_avalon_shell_rsa_0_s0_address;      // mm_interconnect_1:avalon_shell_rsa_0_s0_address -> avalon_shell_rsa_0:avs_s0_address
	wire          mm_interconnect_1_avalon_shell_rsa_0_s0_read;         // mm_interconnect_1:avalon_shell_rsa_0_s0_read -> avalon_shell_rsa_0:avs_s0_read
	wire          mm_interconnect_1_avalon_shell_rsa_0_s0_write;        // mm_interconnect_1:avalon_shell_rsa_0_s0_write -> avalon_shell_rsa_0:avs_s0_write
	wire  [127:0] mm_interconnect_1_avalon_shell_rsa_0_s0_writedata;    // mm_interconnect_1:avalon_shell_rsa_0_s0_writedata -> avalon_shell_rsa_0:avs_s0_writedata
	wire          dma0_pp_m0_waitrequest;                               // mm_interconnect_2:dma0_pp_m0_waitrequest -> dma0_pp:m0_waitrequest
	wire  [127:0] dma0_pp_m0_readdata;                                  // mm_interconnect_2:dma0_pp_m0_readdata -> dma0_pp:m0_readdata
	wire          dma0_pp_m0_debugaccess;                               // dma0_pp:m0_debugaccess -> mm_interconnect_2:dma0_pp_m0_debugaccess
	wire   [31:0] dma0_pp_m0_address;                                   // dma0_pp:m0_address -> mm_interconnect_2:dma0_pp_m0_address
	wire          dma0_pp_m0_read;                                      // dma0_pp:m0_read -> mm_interconnect_2:dma0_pp_m0_read
	wire   [15:0] dma0_pp_m0_byteenable;                                // dma0_pp:m0_byteenable -> mm_interconnect_2:dma0_pp_m0_byteenable
	wire          dma0_pp_m0_readdatavalid;                             // mm_interconnect_2:dma0_pp_m0_readdatavalid -> dma0_pp:m0_readdatavalid
	wire  [127:0] dma0_pp_m0_writedata;                                 // dma0_pp:m0_writedata -> mm_interconnect_2:dma0_pp_m0_writedata
	wire          dma0_pp_m0_write;                                     // dma0_pp:m0_write -> mm_interconnect_2:dma0_pp_m0_write
	wire    [9:0] dma0_pp_m0_burstcount;                                // dma0_pp:m0_burstcount -> mm_interconnect_2:dma0_pp_m0_burstcount
	wire          avalon_shell_rsa_0_m0_waitrequest;                    // mm_interconnect_2:avalon_shell_rsa_0_m0_waitrequest -> avalon_shell_rsa_0:avm_m0_waitrequest
	wire    [7:0] avalon_shell_rsa_0_m0_readdata;                       // mm_interconnect_2:avalon_shell_rsa_0_m0_readdata -> avalon_shell_rsa_0:avm_m0_readdata
	wire   [31:0] avalon_shell_rsa_0_m0_address;                        // avalon_shell_rsa_0:avm_m0_address -> mm_interconnect_2:avalon_shell_rsa_0_m0_address
	wire          avalon_shell_rsa_0_m0_read;                           // avalon_shell_rsa_0:avm_m0_read -> mm_interconnect_2:avalon_shell_rsa_0_m0_read
	wire          avalon_shell_rsa_0_m0_write;                          // avalon_shell_rsa_0:avm_m0_write -> mm_interconnect_2:avalon_shell_rsa_0_m0_write
	wire    [7:0] avalon_shell_rsa_0_m0_writedata;                      // avalon_shell_rsa_0:avm_m0_writedata -> mm_interconnect_2:avalon_shell_rsa_0_m0_writedata
	wire          mm_interconnect_2_pcie_interface_txs_chipselect;      // mm_interconnect_2:PCIE_interface_Txs_chipselect -> PCIE_interface:TxsChipSelect_i
	wire  [127:0] mm_interconnect_2_pcie_interface_txs_readdata;        // PCIE_interface:TxsReadData_o -> mm_interconnect_2:PCIE_interface_Txs_readdata
	wire          mm_interconnect_2_pcie_interface_txs_waitrequest;     // PCIE_interface:TxsWaitRequest_o -> mm_interconnect_2:PCIE_interface_Txs_waitrequest
	wire   [30:0] mm_interconnect_2_pcie_interface_txs_address;         // mm_interconnect_2:PCIE_interface_Txs_address -> PCIE_interface:TxsAddress_i
	wire          mm_interconnect_2_pcie_interface_txs_read;            // mm_interconnect_2:PCIE_interface_Txs_read -> PCIE_interface:TxsRead_i
	wire   [15:0] mm_interconnect_2_pcie_interface_txs_byteenable;      // mm_interconnect_2:PCIE_interface_Txs_byteenable -> PCIE_interface:TxsByteEnable_i
	wire          mm_interconnect_2_pcie_interface_txs_readdatavalid;   // PCIE_interface:TxsReadDataValid_o -> mm_interconnect_2:PCIE_interface_Txs_readdatavalid
	wire          mm_interconnect_2_pcie_interface_txs_write;           // mm_interconnect_2:PCIE_interface_Txs_write -> PCIE_interface:TxsWrite_i
	wire  [127:0] mm_interconnect_2_pcie_interface_txs_writedata;       // mm_interconnect_2:PCIE_interface_Txs_writedata -> PCIE_interface:TxsWriteData_i
	wire    [5:0] mm_interconnect_2_pcie_interface_txs_burstcount;      // mm_interconnect_2:PCIE_interface_Txs_burstcount -> PCIE_interface:TxsBurstCount_i
	wire          mm_interconnect_2_ddr3a_avl_beginbursttransfer;       // mm_interconnect_2:ddr3a_avl_beginbursttransfer -> ddr3a:avl_burstbegin
	wire  [511:0] mm_interconnect_2_ddr3a_avl_readdata;                 // ddr3a:avl_rdata -> mm_interconnect_2:ddr3a_avl_readdata
	wire          mm_interconnect_2_ddr3a_avl_waitrequest;              // ddr3a:avl_ready -> mm_interconnect_2:ddr3a_avl_waitrequest
	wire   [24:0] mm_interconnect_2_ddr3a_avl_address;                  // mm_interconnect_2:ddr3a_avl_address -> ddr3a:avl_addr
	wire          mm_interconnect_2_ddr3a_avl_read;                     // mm_interconnect_2:ddr3a_avl_read -> ddr3a:avl_read_req
	wire   [63:0] mm_interconnect_2_ddr3a_avl_byteenable;               // mm_interconnect_2:ddr3a_avl_byteenable -> ddr3a:avl_be
	wire          mm_interconnect_2_ddr3a_avl_readdatavalid;            // ddr3a:avl_rdata_valid -> mm_interconnect_2:ddr3a_avl_readdatavalid
	wire          mm_interconnect_2_ddr3a_avl_write;                    // mm_interconnect_2:ddr3a_avl_write -> ddr3a:avl_write_req
	wire  [511:0] mm_interconnect_2_ddr3a_avl_writedata;                // mm_interconnect_2:ddr3a_avl_writedata -> ddr3a:avl_wdata
	wire    [9:0] mm_interconnect_2_ddr3a_avl_burstcount;               // mm_interconnect_2:ddr3a_avl_burstcount -> ddr3a:avl_size
	wire          ddr3a_afi_clk_clk;                                    // ddr3a:afi_clk -> [mm_interconnect_2:ddr3a_afi_clk_clk, rst_controller_002:clk]
	wire          dma0_read_master_chipselect;                          // dma0:read_chipselect -> mm_interconnect_3:dma0_read_master_chipselect
	wire  [127:0] dma0_read_master_readdata;                            // mm_interconnect_3:dma0_read_master_readdata -> dma0:read_readdata
	wire          dma0_read_master_waitrequest;                         // mm_interconnect_3:dma0_read_master_waitrequest -> dma0:read_waitrequest
	wire   [31:0] dma0_read_master_address;                             // dma0:read_address -> mm_interconnect_3:dma0_read_master_address
	wire          dma0_read_master_read;                                // dma0:read_read_n -> mm_interconnect_3:dma0_read_master_read
	wire          dma0_read_master_readdatavalid;                       // mm_interconnect_3:dma0_read_master_readdatavalid -> dma0:read_readdatavalid
	wire    [9:0] dma0_read_master_burstcount;                          // dma0:read_burstcount -> mm_interconnect_3:dma0_read_master_burstcount
	wire          dma0_write_master_chipselect;                         // dma0:write_chipselect -> mm_interconnect_3:dma0_write_master_chipselect
	wire          dma0_write_master_waitrequest;                        // mm_interconnect_3:dma0_write_master_waitrequest -> dma0:write_waitrequest
	wire   [31:0] dma0_write_master_address;                            // dma0:write_address -> mm_interconnect_3:dma0_write_master_address
	wire   [15:0] dma0_write_master_byteenable;                         // dma0:write_byteenable -> mm_interconnect_3:dma0_write_master_byteenable
	wire          dma0_write_master_write;                              // dma0:write_write_n -> mm_interconnect_3:dma0_write_master_write
	wire  [127:0] dma0_write_master_writedata;                          // dma0:write_writedata -> mm_interconnect_3:dma0_write_master_writedata
	wire    [9:0] dma0_write_master_burstcount;                         // dma0:write_burstcount -> mm_interconnect_3:dma0_write_master_burstcount
	wire  [127:0] mm_interconnect_3_dma0_pp_s0_readdata;                // dma0_pp:s0_readdata -> mm_interconnect_3:dma0_pp_s0_readdata
	wire          mm_interconnect_3_dma0_pp_s0_waitrequest;             // dma0_pp:s0_waitrequest -> mm_interconnect_3:dma0_pp_s0_waitrequest
	wire          mm_interconnect_3_dma0_pp_s0_debugaccess;             // mm_interconnect_3:dma0_pp_s0_debugaccess -> dma0_pp:s0_debugaccess
	wire   [31:0] mm_interconnect_3_dma0_pp_s0_address;                 // mm_interconnect_3:dma0_pp_s0_address -> dma0_pp:s0_address
	wire          mm_interconnect_3_dma0_pp_s0_read;                    // mm_interconnect_3:dma0_pp_s0_read -> dma0_pp:s0_read
	wire   [15:0] mm_interconnect_3_dma0_pp_s0_byteenable;              // mm_interconnect_3:dma0_pp_s0_byteenable -> dma0_pp:s0_byteenable
	wire          mm_interconnect_3_dma0_pp_s0_readdatavalid;           // dma0_pp:s0_readdatavalid -> mm_interconnect_3:dma0_pp_s0_readdatavalid
	wire          mm_interconnect_3_dma0_pp_s0_write;                   // mm_interconnect_3:dma0_pp_s0_write -> dma0_pp:s0_write
	wire  [127:0] mm_interconnect_3_dma0_pp_s0_writedata;               // mm_interconnect_3:dma0_pp_s0_writedata -> dma0_pp:s0_writedata
	wire    [9:0] mm_interconnect_3_dma0_pp_s0_burstcount;              // mm_interconnect_3:dma0_pp_s0_burstcount -> dma0_pp:s0_burstcount
	wire          irq_mapper_receiver0_irq;                             // dma0:dma_ctl_irq -> irq_mapper:receiver0_irq
	wire   [15:0] pcie_interface_rxmirq_irq;                            // irq_mapper:sender_irq -> PCIE_interface:RxmIrq_i
	wire          rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [PCIe_config:mgmt_rst_reset, PCIe_config_driver:reconfig_xcvr_rst, avalon_shell_rsa_0:reset, mm_interconnect_1:avalon_shell_rsa_0_reset_reset_bridge_in_reset_reset, mm_interconnect_2:avalon_shell_rsa_0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                   // rst_controller_001:reset_out -> [dma0:system_reset_n, dma0_pp:reset, irq_mapper:reset, mm_interconnect_0:dma0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:PCIE_interface_Rxm_BAR2_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:dma0_pp_reset_reset_bridge_in_reset_reset, mm_interconnect_3:dma0_reset_reset_bridge_in_reset_reset]
	wire          pcie_interface_nreset_status_reset;                   // PCIE_interface:reset_status -> rst_controller_001:reset_in0
	wire          rst_controller_002_reset_out_reset;                   // rst_controller_002:reset_out -> [mm_interconnect_2:ddr3a_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_2:ddr3a_soft_reset_reset_bridge_in_reset_reset]

	altpcie_sv_hip_avmm_hwtcl #(
		.lane_mask_hwtcl                          ("x8"),
		.gen123_lane_rate_mode_hwtcl              ("Gen2 (5.0 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("2.1"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.in_cvp_mode_hwtcl                        (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.use_atx_pll_hwtcl                        (0),
		.enable_power_on_rst_pulse_hwtcl          (0),
		.enable_pcisigtest_hwtcl                  (0),
		.bar0_size_mask_hwtcl                     (15),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Disabled"),
		.bar0_prefetchable_hwtcl                  ("Disabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (5),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Disabled"),
		.bar2_prefetchable_hwtcl                  ("Disabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (0),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Disabled"),
		.bar4_prefetchable_hwtcl                  ("Disabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.vendor_id_hwtcl                          (4466),
		.device_id_hwtcl                          (21862),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (0),
		.subsystem_vendor_id_hwtcl                (9509),
		.subsystem_device_id_hwtcl                (9509),
		.max_payload_size_hwtcl                   (256),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (0),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.avmm_width_hwtcl                         (128),
		.AVALON_ADDR_WIDTH                        (32),
		.avmm_burst_width_hwtcl                   (6),
		.CB_PCIE_MODE                             (0),
		.CB_PCIE_RX_LITE                          (0),
		.CB_RXM_DATA_WIDTH                        (128),
		.CG_AVALON_S_ADDR_WIDTH                   (31),
		.CG_IMPL_CRA_AV_SLAVE_PORT                (1),
		.CG_ENABLE_ADVANCED_INTERRUPT             (0),
		.CG_ENABLE_A2P_INTERRUPT                  (0),
		.CB_A2P_ADDR_MAP_IS_FIXED                 (0),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES              (2),
		.BYPASSS_A2P_TRANSLATION                  (0),
		.a2p_pass_thru_bits                       (30),
		.ast_width_hwtcl                          ("Avalon-ST 128-bit"),
		.use_ast_parity                           (0),
		.millisecond_cycle_count_hwtcl            (248500),
		.port_width_be_hwtcl                      (16),
		.port_width_data_hwtcl                    (128),
		.hip_reconfig_hwtcl                       (0),
		.vsec_id_hwtcl                            (40960),
		.vsec_rev_hwtcl                           (0),
		.expansion_base_address_register_hwtcl    (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("true"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (195),
		.cpl_spc_data_hwtcl                       (781),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("config_retry_status"),
		.core_clk_sel_hwtcl                       ("pld_clk"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (700),
		.reconfig_from_xcvr_width                 (460),
		.single_rx_detect_hwtcl                   (0),
		.hip_hard_reset_hwtcl                     (0),
		.use_cvp_update_core_pof_hwtcl            (0),
		.pcie_inspector_hwtcl                     (0),
		.tlp_inspector_hwtcl                      (0),
		.tlp_inspector_use_signal_probe_hwtcl     (0),
		.tlp_insp_trg_dw0_hwtcl                   (2049),
		.tlp_insp_trg_dw1_hwtcl                   (0),
		.tlp_insp_trg_dw2_hwtcl                   (0),
		.tlp_insp_trg_dw3_hwtcl                   (0),
		.hwtcl_override_g2_txvod                  (1),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15)
	) pcie_interface (
		.coreclkout           (pcie_interface_coreclkout_clk),                        //          coreclkout.clk
		.refclk               (pcie_interface_refclk_clk),                            //              refclk.clk
		.npor                 (pcie_interface_npor_npor),                             //                npor.npor
		.pin_perst            (pcie_interface_npor_pin_perst),                        //                    .pin_perst
		.reset_status         (pcie_interface_nreset_status_reset),                   //       nreset_status.reset_n
		.RxmAddress_0_o       (pcie_interface_rxm_bar0_address),                      //            Rxm_BAR0.address
		.RxmRead_0_o          (pcie_interface_rxm_bar0_read),                         //                    .read
		.RxmWaitRequest_0_i   (pcie_interface_rxm_bar0_waitrequest),                  //                    .waitrequest
		.RxmWrite_0_o         (pcie_interface_rxm_bar0_write),                        //                    .write
		.RxmReadDataValid_0_i (pcie_interface_rxm_bar0_readdatavalid),                //                    .readdatavalid
		.RxmReadData_0_i      (pcie_interface_rxm_bar0_readdata),                     //                    .readdata
		.RxmWriteData_0_o     (pcie_interface_rxm_bar0_writedata),                    //                    .writedata
		.RxmBurstCount_0_o    (pcie_interface_rxm_bar0_burstcount),                   //                    .burstcount
		.RxmByteEnable_0_o    (pcie_interface_rxm_bar0_byteenable),                   //                    .byteenable
		.RxmAddress_2_o       (pcie_interface_rxm_bar2_address),                      //            Rxm_BAR2.address
		.RxmRead_2_o          (pcie_interface_rxm_bar2_read),                         //                    .read
		.RxmWaitRequest_2_i   (pcie_interface_rxm_bar2_waitrequest),                  //                    .waitrequest
		.RxmWrite_2_o         (pcie_interface_rxm_bar2_write),                        //                    .write
		.RxmReadDataValid_2_i (pcie_interface_rxm_bar2_readdatavalid),                //                    .readdatavalid
		.RxmReadData_2_i      (pcie_interface_rxm_bar2_readdata),                     //                    .readdata
		.RxmWriteData_2_o     (pcie_interface_rxm_bar2_writedata),                    //                    .writedata
		.RxmBurstCount_2_o    (pcie_interface_rxm_bar2_burstcount),                   //                    .burstcount
		.RxmByteEnable_2_o    (pcie_interface_rxm_bar2_byteenable),                   //                    .byteenable
		.RxmIrq_i             (pcie_interface_rxmirq_irq),                            //              RxmIrq.irq
		.derr_cor_ext_rcv     (pcie_interface_hip_status_derr_cor_ext_rcv),           //          hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl     (pcie_interface_hip_status_derr_cor_ext_rpl),           //                    .derr_cor_ext_rpl
		.derr_rpl             (pcie_interface_hip_status_derr_rpl),                   //                    .derr_rpl
		.dlup                 (pcie_interface_hip_status_dlup),                       //                    .dlup
		.dlup_exit            (pcie_interface_hip_status_dlup_exit),                  //                    .dlup_exit
		.ev128ns              (pcie_interface_hip_status_ev128ns),                    //                    .ev128ns
		.ev1us                (pcie_interface_hip_status_ev1us),                      //                    .ev1us
		.hotrst_exit          (pcie_interface_hip_status_hotrst_exit),                //                    .hotrst_exit
		.int_status           (pcie_interface_hip_status_int_status),                 //                    .int_status
		.l2_exit              (pcie_interface_hip_status_l2_exit),                    //                    .l2_exit
		.lane_act             (pcie_interface_hip_status_lane_act),                   //                    .lane_act
		.ltssmstate           (pcie_interface_hip_status_ltssmstate),                 //                    .ltssmstate
		.rx_par_err           (pcie_interface_hip_status_rx_par_err),                 //                    .rx_par_err
		.tx_par_err           (pcie_interface_hip_status_tx_par_err),                 //                    .tx_par_err
		.cfg_par_err          (pcie_interface_hip_status_cfg_par_err),                //                    .cfg_par_err
		.ko_cpl_spc_header    (pcie_interface_hip_status_ko_cpl_spc_header),          //                    .ko_cpl_spc_header
		.ko_cpl_spc_data      (pcie_interface_hip_status_ko_cpl_spc_data),            //                    .ko_cpl_spc_data
		.currentspeed         (pcie_interface_hip_currentspeed_currentspeed),         //    hip_currentspeed.currentspeed
		.reconfig_to_xcvr     (pcie_config_reconfig_to_xcvr_reconfig_to_xcvr),        //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr   (pcie_interface_reconfig_from_xcvr_reconfig_from_xcvr), //  reconfig_from_xcvr.reconfig_from_xcvr
		.fixedclk_locked      (),                                                     // reconfig_clk_locked.fixedclk_locked
		.rx_in0               (pcie_interface_hip_serial_rx_in0),                     //          hip_serial.rx_in0
		.rx_in1               (pcie_interface_hip_serial_rx_in1),                     //                    .rx_in1
		.rx_in2               (pcie_interface_hip_serial_rx_in2),                     //                    .rx_in2
		.rx_in3               (pcie_interface_hip_serial_rx_in3),                     //                    .rx_in3
		.rx_in4               (pcie_interface_hip_serial_rx_in4),                     //                    .rx_in4
		.rx_in5               (pcie_interface_hip_serial_rx_in5),                     //                    .rx_in5
		.rx_in6               (pcie_interface_hip_serial_rx_in6),                     //                    .rx_in6
		.rx_in7               (pcie_interface_hip_serial_rx_in7),                     //                    .rx_in7
		.tx_out0              (pcie_interface_hip_serial_tx_out0),                    //                    .tx_out0
		.tx_out1              (pcie_interface_hip_serial_tx_out1),                    //                    .tx_out1
		.tx_out2              (pcie_interface_hip_serial_tx_out2),                    //                    .tx_out2
		.tx_out3              (pcie_interface_hip_serial_tx_out3),                    //                    .tx_out3
		.tx_out4              (pcie_interface_hip_serial_tx_out4),                    //                    .tx_out4
		.tx_out5              (pcie_interface_hip_serial_tx_out5),                    //                    .tx_out5
		.tx_out6              (pcie_interface_hip_serial_tx_out6),                    //                    .tx_out6
		.tx_out7              (pcie_interface_hip_serial_tx_out7),                    //                    .tx_out7
		.sim_pipe_pclk_in     (),                                                     //            hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate        (),                                                     //                    .sim_pipe_rate
		.sim_ltssmstate       (),                                                     //                    .sim_ltssmstate
		.eidleinfersel0       (),                                                     //                    .eidleinfersel0
		.eidleinfersel1       (),                                                     //                    .eidleinfersel1
		.eidleinfersel2       (),                                                     //                    .eidleinfersel2
		.eidleinfersel3       (),                                                     //                    .eidleinfersel3
		.eidleinfersel4       (),                                                     //                    .eidleinfersel4
		.eidleinfersel5       (),                                                     //                    .eidleinfersel5
		.eidleinfersel6       (),                                                     //                    .eidleinfersel6
		.eidleinfersel7       (),                                                     //                    .eidleinfersel7
		.powerdown0           (),                                                     //                    .powerdown0
		.powerdown1           (),                                                     //                    .powerdown1
		.powerdown2           (),                                                     //                    .powerdown2
		.powerdown3           (),                                                     //                    .powerdown3
		.powerdown4           (),                                                     //                    .powerdown4
		.powerdown5           (),                                                     //                    .powerdown5
		.powerdown6           (),                                                     //                    .powerdown6
		.powerdown7           (),                                                     //                    .powerdown7
		.rxpolarity0          (),                                                     //                    .rxpolarity0
		.rxpolarity1          (),                                                     //                    .rxpolarity1
		.rxpolarity2          (),                                                     //                    .rxpolarity2
		.rxpolarity3          (),                                                     //                    .rxpolarity3
		.rxpolarity4          (),                                                     //                    .rxpolarity4
		.rxpolarity5          (),                                                     //                    .rxpolarity5
		.rxpolarity6          (),                                                     //                    .rxpolarity6
		.rxpolarity7          (),                                                     //                    .rxpolarity7
		.txcompl0             (),                                                     //                    .txcompl0
		.txcompl1             (),                                                     //                    .txcompl1
		.txcompl2             (),                                                     //                    .txcompl2
		.txcompl3             (),                                                     //                    .txcompl3
		.txcompl4             (),                                                     //                    .txcompl4
		.txcompl5             (),                                                     //                    .txcompl5
		.txcompl6             (),                                                     //                    .txcompl6
		.txcompl7             (),                                                     //                    .txcompl7
		.txdata0              (),                                                     //                    .txdata0
		.txdata1              (),                                                     //                    .txdata1
		.txdata2              (),                                                     //                    .txdata2
		.txdata3              (),                                                     //                    .txdata3
		.txdata4              (),                                                     //                    .txdata4
		.txdata5              (),                                                     //                    .txdata5
		.txdata6              (),                                                     //                    .txdata6
		.txdata7              (),                                                     //                    .txdata7
		.txdatak0             (),                                                     //                    .txdatak0
		.txdatak1             (),                                                     //                    .txdatak1
		.txdatak2             (),                                                     //                    .txdatak2
		.txdatak3             (),                                                     //                    .txdatak3
		.txdatak4             (),                                                     //                    .txdatak4
		.txdatak5             (),                                                     //                    .txdatak5
		.txdatak6             (),                                                     //                    .txdatak6
		.txdatak7             (),                                                     //                    .txdatak7
		.txdetectrx0          (),                                                     //                    .txdetectrx0
		.txdetectrx1          (),                                                     //                    .txdetectrx1
		.txdetectrx2          (),                                                     //                    .txdetectrx2
		.txdetectrx3          (),                                                     //                    .txdetectrx3
		.txdetectrx4          (),                                                     //                    .txdetectrx4
		.txdetectrx5          (),                                                     //                    .txdetectrx5
		.txdetectrx6          (),                                                     //                    .txdetectrx6
		.txdetectrx7          (),                                                     //                    .txdetectrx7
		.txelecidle0          (),                                                     //                    .txelecidle0
		.txelecidle1          (),                                                     //                    .txelecidle1
		.txelecidle2          (),                                                     //                    .txelecidle2
		.txelecidle3          (),                                                     //                    .txelecidle3
		.txelecidle4          (),                                                     //                    .txelecidle4
		.txelecidle5          (),                                                     //                    .txelecidle5
		.txelecidle6          (),                                                     //                    .txelecidle6
		.txelecidle7          (),                                                     //                    .txelecidle7
		.txdeemph0            (),                                                     //                    .txdeemph0
		.txdeemph1            (),                                                     //                    .txdeemph1
		.txdeemph2            (),                                                     //                    .txdeemph2
		.txdeemph3            (),                                                     //                    .txdeemph3
		.txdeemph4            (),                                                     //                    .txdeemph4
		.txdeemph5            (),                                                     //                    .txdeemph5
		.txdeemph6            (),                                                     //                    .txdeemph6
		.txdeemph7            (),                                                     //                    .txdeemph7
		.txmargin0            (),                                                     //                    .txmargin0
		.txmargin1            (),                                                     //                    .txmargin1
		.txmargin2            (),                                                     //                    .txmargin2
		.txmargin3            (),                                                     //                    .txmargin3
		.txmargin4            (),                                                     //                    .txmargin4
		.txmargin5            (),                                                     //                    .txmargin5
		.txmargin6            (),                                                     //                    .txmargin6
		.txmargin7            (),                                                     //                    .txmargin7
		.txswing0             (),                                                     //                    .txswing0
		.txswing1             (),                                                     //                    .txswing1
		.txswing2             (),                                                     //                    .txswing2
		.txswing3             (),                                                     //                    .txswing3
		.txswing4             (),                                                     //                    .txswing4
		.txswing5             (),                                                     //                    .txswing5
		.txswing6             (),                                                     //                    .txswing6
		.txswing7             (),                                                     //                    .txswing7
		.phystatus0           (),                                                     //                    .phystatus0
		.phystatus1           (),                                                     //                    .phystatus1
		.phystatus2           (),                                                     //                    .phystatus2
		.phystatus3           (),                                                     //                    .phystatus3
		.phystatus4           (),                                                     //                    .phystatus4
		.phystatus5           (),                                                     //                    .phystatus5
		.phystatus6           (),                                                     //                    .phystatus6
		.phystatus7           (),                                                     //                    .phystatus7
		.rxdata0              (),                                                     //                    .rxdata0
		.rxdata1              (),                                                     //                    .rxdata1
		.rxdata2              (),                                                     //                    .rxdata2
		.rxdata3              (),                                                     //                    .rxdata3
		.rxdata4              (),                                                     //                    .rxdata4
		.rxdata5              (),                                                     //                    .rxdata5
		.rxdata6              (),                                                     //                    .rxdata6
		.rxdata7              (),                                                     //                    .rxdata7
		.rxdatak0             (),                                                     //                    .rxdatak0
		.rxdatak1             (),                                                     //                    .rxdatak1
		.rxdatak2             (),                                                     //                    .rxdatak2
		.rxdatak3             (),                                                     //                    .rxdatak3
		.rxdatak4             (),                                                     //                    .rxdatak4
		.rxdatak5             (),                                                     //                    .rxdatak5
		.rxdatak6             (),                                                     //                    .rxdatak6
		.rxdatak7             (),                                                     //                    .rxdatak7
		.rxelecidle0          (),                                                     //                    .rxelecidle0
		.rxelecidle1          (),                                                     //                    .rxelecidle1
		.rxelecidle2          (),                                                     //                    .rxelecidle2
		.rxelecidle3          (),                                                     //                    .rxelecidle3
		.rxelecidle4          (),                                                     //                    .rxelecidle4
		.rxelecidle5          (),                                                     //                    .rxelecidle5
		.rxelecidle6          (),                                                     //                    .rxelecidle6
		.rxelecidle7          (),                                                     //                    .rxelecidle7
		.rxstatus0            (),                                                     //                    .rxstatus0
		.rxstatus1            (),                                                     //                    .rxstatus1
		.rxstatus2            (),                                                     //                    .rxstatus2
		.rxstatus3            (),                                                     //                    .rxstatus3
		.rxstatus4            (),                                                     //                    .rxstatus4
		.rxstatus5            (),                                                     //                    .rxstatus5
		.rxstatus6            (),                                                     //                    .rxstatus6
		.rxstatus7            (),                                                     //                    .rxstatus7
		.rxvalid0             (),                                                     //                    .rxvalid0
		.rxvalid1             (),                                                     //                    .rxvalid1
		.rxvalid2             (),                                                     //                    .rxvalid2
		.rxvalid3             (),                                                     //                    .rxvalid3
		.rxvalid4             (),                                                     //                    .rxvalid4
		.rxvalid5             (),                                                     //                    .rxvalid5
		.rxvalid6             (),                                                     //                    .rxvalid6
		.rxvalid7             (),                                                     //                    .rxvalid7
		.test_in              (),                                                     //            hip_ctrl.test_in
		.simu_mode_pipe       (),                                                     //                    .simu_mode_pipe
		.TxsChipSelect_i      (mm_interconnect_2_pcie_interface_txs_chipselect),      //                 Txs.chipselect
		.TxsByteEnable_i      (mm_interconnect_2_pcie_interface_txs_byteenable),      //                    .byteenable
		.TxsReadData_o        (mm_interconnect_2_pcie_interface_txs_readdata),        //                    .readdata
		.TxsWriteData_i       (mm_interconnect_2_pcie_interface_txs_writedata),       //                    .writedata
		.TxsRead_i            (mm_interconnect_2_pcie_interface_txs_read),            //                    .read
		.TxsWrite_i           (mm_interconnect_2_pcie_interface_txs_write),           //                    .write
		.TxsBurstCount_i      (mm_interconnect_2_pcie_interface_txs_burstcount),      //                    .burstcount
		.TxsReadDataValid_o   (mm_interconnect_2_pcie_interface_txs_readdatavalid),   //                    .readdatavalid
		.TxsWaitRequest_o     (mm_interconnect_2_pcie_interface_txs_waitrequest),     //                    .waitrequest
		.TxsAddress_i         (mm_interconnect_2_pcie_interface_txs_address),         //                    .address
		.CraChipSelect_i      (mm_interconnect_0_pcie_interface_cra_chipselect),      //                 Cra.chipselect
		.CraAddress_i         (mm_interconnect_0_pcie_interface_cra_address),         //                    .address
		.CraByteEnable_i      (mm_interconnect_0_pcie_interface_cra_byteenable),      //                    .byteenable
		.CraRead              (mm_interconnect_0_pcie_interface_cra_read),            //                    .read
		.CraReadData_o        (mm_interconnect_0_pcie_interface_cra_readdata),        //                    .readdata
		.CraWrite             (mm_interconnect_0_pcie_interface_cra_write),           //                    .write
		.CraWriteData_i       (mm_interconnect_0_pcie_interface_cra_writedata),       //                    .writedata
		.CraWaitRequest_o     (mm_interconnect_0_pcie_interface_cra_waitrequest),     //                    .waitrequest
		.CraIrq_o             (),                                                     //              CraIrq.irq
		.rxdataskip0          (1'b0),                                                 //         (terminated)
		.rxdataskip1          (1'b0),                                                 //         (terminated)
		.rxdataskip2          (1'b0),                                                 //         (terminated)
		.rxdataskip3          (1'b0),                                                 //         (terminated)
		.rxdataskip4          (1'b0),                                                 //         (terminated)
		.rxdataskip5          (1'b0),                                                 //         (terminated)
		.rxdataskip6          (1'b0),                                                 //         (terminated)
		.rxdataskip7          (1'b0),                                                 //         (terminated)
		.rxblkst0             (1'b0),                                                 //         (terminated)
		.rxblkst1             (1'b0),                                                 //         (terminated)
		.rxblkst2             (1'b0),                                                 //         (terminated)
		.rxblkst3             (1'b0),                                                 //         (terminated)
		.rxblkst4             (1'b0),                                                 //         (terminated)
		.rxblkst5             (1'b0),                                                 //         (terminated)
		.rxblkst6             (1'b0),                                                 //         (terminated)
		.rxblkst7             (1'b0),                                                 //         (terminated)
		.rxsynchd0            (2'b00),                                                //         (terminated)
		.rxsynchd1            (2'b00),                                                //         (terminated)
		.rxsynchd2            (2'b00),                                                //         (terminated)
		.rxsynchd3            (2'b00),                                                //         (terminated)
		.rxsynchd4            (2'b00),                                                //         (terminated)
		.rxsynchd5            (2'b00),                                                //         (terminated)
		.rxsynchd6            (2'b00),                                                //         (terminated)
		.rxsynchd7            (2'b00),                                                //         (terminated)
		.rxfreqlocked0        (1'b0),                                                 //         (terminated)
		.rxfreqlocked1        (1'b0),                                                 //         (terminated)
		.rxfreqlocked2        (1'b0),                                                 //         (terminated)
		.rxfreqlocked3        (1'b0),                                                 //         (terminated)
		.rxfreqlocked4        (1'b0),                                                 //         (terminated)
		.rxfreqlocked5        (1'b0),                                                 //         (terminated)
		.rxfreqlocked6        (1'b0),                                                 //         (terminated)
		.rxfreqlocked7        (1'b0),                                                 //         (terminated)
		.currentcoeff0        (),                                                     //         (terminated)
		.currentcoeff1        (),                                                     //         (terminated)
		.currentcoeff2        (),                                                     //         (terminated)
		.currentcoeff3        (),                                                     //         (terminated)
		.currentcoeff4        (),                                                     //         (terminated)
		.currentcoeff5        (),                                                     //         (terminated)
		.currentcoeff6        (),                                                     //         (terminated)
		.currentcoeff7        (),                                                     //         (terminated)
		.currentrxpreset0     (),                                                     //         (terminated)
		.currentrxpreset1     (),                                                     //         (terminated)
		.currentrxpreset2     (),                                                     //         (terminated)
		.currentrxpreset3     (),                                                     //         (terminated)
		.currentrxpreset4     (),                                                     //         (terminated)
		.currentrxpreset5     (),                                                     //         (terminated)
		.currentrxpreset6     (),                                                     //         (terminated)
		.currentrxpreset7     (),                                                     //         (terminated)
		.txsynchd0            (),                                                     //         (terminated)
		.txsynchd1            (),                                                     //         (terminated)
		.txsynchd2            (),                                                     //         (terminated)
		.txsynchd3            (),                                                     //         (terminated)
		.txsynchd4            (),                                                     //         (terminated)
		.txsynchd5            (),                                                     //         (terminated)
		.txsynchd6            (),                                                     //         (terminated)
		.txsynchd7            (),                                                     //         (terminated)
		.txblkst0             (),                                                     //         (terminated)
		.txblkst1             (),                                                     //         (terminated)
		.txblkst2             (),                                                     //         (terminated)
		.txblkst3             (),                                                     //         (terminated)
		.txblkst4             (),                                                     //         (terminated)
		.txblkst5             (),                                                     //         (terminated)
		.txblkst6             (),                                                     //         (terminated)
		.txblkst7             ()                                                      //         (terminated)
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (10),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (1),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) pcie_config (
		.reconfig_busy             (pcie_config_reconfig_busy_reconfig_busy),              //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_0_clk),                                            //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_reset_out_reset),                       //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (pcie_config_driver_reconfig_mgmt_address),             //      reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_config_driver_reconfig_mgmt_read),                //                   .read
		.reconfig_mgmt_readdata    (pcie_config_driver_reconfig_mgmt_readdata),            //                   .readdata
		.reconfig_mgmt_waitrequest (pcie_config_driver_reconfig_mgmt_waitrequest),         //                   .waitrequest
		.reconfig_mgmt_write       (pcie_config_driver_reconfig_mgmt_write),               //                   .write
		.reconfig_mgmt_writedata   (pcie_config_driver_reconfig_mgmt_writedata),           //                   .writedata
		.reconfig_to_xcvr          (pcie_config_reconfig_to_xcvr_reconfig_to_xcvr),        //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (pcie_interface_reconfig_from_xcvr_reconfig_from_xcvr), // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                     //        (terminated)
		.rx_cal_busy               (),                                                     //        (terminated)
		.cal_busy_in               (1'b0),                                                 //        (terminated)
		.reconfig_mif_address      (),                                                     //        (terminated)
		.reconfig_mif_read         (),                                                     //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                                 //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                                  //        (terminated)
	);

	altpcie_reconfig_driver #(
		.INTENDED_DEVICE_FAMILY        ("Stratix V"),
		.gen123_lane_rate_mode_hwtcl   ("Gen2 (5.0 Gbps)"),
		.number_of_reconfig_interfaces (10)
	) pcie_config_driver (
		.reconfig_xcvr_clk         (clk_0_clk),                                    // reconfig_xcvr_clk.clk
		.reconfig_xcvr_rst         (rst_controller_reset_out_reset),               // reconfig_xcvr_rst.reset
		.reconfig_mgmt_address     (pcie_config_driver_reconfig_mgmt_address),     //     reconfig_mgmt.address
		.reconfig_mgmt_read        (pcie_config_driver_reconfig_mgmt_read),        //                  .read
		.reconfig_mgmt_readdata    (pcie_config_driver_reconfig_mgmt_readdata),    //                  .readdata
		.reconfig_mgmt_waitrequest (pcie_config_driver_reconfig_mgmt_waitrequest), //                  .waitrequest
		.reconfig_mgmt_write       (pcie_config_driver_reconfig_mgmt_write),       //                  .write
		.reconfig_mgmt_writedata   (pcie_config_driver_reconfig_mgmt_writedata),   //                  .writedata
		.currentspeed              (pcie_interface_hip_currentspeed_currentspeed), //  hip_currentspeed.currentspeed
		.reconfig_busy             (pcie_config_reconfig_busy_reconfig_busy),      //     reconfig_busy.reconfig_busy
		.pld_clk                   (pcie_interface_coreclkout_clk),                //           pld_clk.clk
		.derr_cor_ext_rcv_drv      (pcie_interface_hip_status_derr_cor_ext_rcv),   //    hip_status_drv.derr_cor_ext_rcv
		.derr_cor_ext_rpl_drv      (pcie_interface_hip_status_derr_cor_ext_rpl),   //                  .derr_cor_ext_rpl
		.derr_rpl_drv              (pcie_interface_hip_status_derr_rpl),           //                  .derr_rpl
		.dlup_exit_drv             (pcie_interface_hip_status_dlup_exit),          //                  .dlup_exit
		.ev128ns_drv               (pcie_interface_hip_status_ev128ns),            //                  .ev128ns
		.ev1us_drv                 (pcie_interface_hip_status_ev1us),              //                  .ev1us
		.hotrst_exit_drv           (pcie_interface_hip_status_hotrst_exit),        //                  .hotrst_exit
		.int_status_drv            (pcie_interface_hip_status_int_status),         //                  .int_status
		.l2_exit_drv               (pcie_interface_hip_status_l2_exit),            //                  .l2_exit
		.lane_act_drv              (pcie_interface_hip_status_lane_act),           //                  .lane_act
		.ltssmstate_drv            (pcie_interface_hip_status_ltssmstate),         //                  .ltssmstate
		.dlup_drv                  (pcie_interface_hip_status_dlup),               //                  .dlup
		.rx_par_err_drv            (pcie_interface_hip_status_rx_par_err),         //                  .rx_par_err
		.tx_par_err_drv            (pcie_interface_hip_status_tx_par_err),         //                  .tx_par_err
		.cfg_par_err_drv           (pcie_interface_hip_status_cfg_par_err),        //                  .cfg_par_err
		.ko_cpl_spc_header_drv     (pcie_interface_hip_status_ko_cpl_spc_header),  //                  .ko_cpl_spc_header
		.ko_cpl_spc_data_drv       (pcie_interface_hip_status_ko_cpl_spc_data),    //                  .ko_cpl_spc_data
		.cal_busy_in               ()                                              //       (terminated)
	);

	avalon_shell_rsa avalon_shell_rsa_0 (
		.clk                       (clk_0_clk),                                           //          clock.clk
		.reset                     (rst_controller_reset_out_reset),                      //          reset.reset
		.avm_m0_waitrequest        (avalon_shell_rsa_0_m0_waitrequest),                   //             m0.waitrequest
		.avm_m0_address            (avalon_shell_rsa_0_m0_address),                       //               .address
		.avm_m0_read               (avalon_shell_rsa_0_m0_read),                          //               .read
		.avm_m0_write              (avalon_shell_rsa_0_m0_write),                         //               .write
		.avm_m0_readdata           (avalon_shell_rsa_0_m0_readdata),                      //               .readdata
		.avm_m0_writedata          (avalon_shell_rsa_0_m0_writedata),                     //               .writedata
		.avs_s0_waitrequest        (mm_interconnect_1_avalon_shell_rsa_0_s0_waitrequest), //             s0.waitrequest
		.avs_s0_address            (mm_interconnect_1_avalon_shell_rsa_0_s0_address),     //               .address
		.avs_s0_read               (mm_interconnect_1_avalon_shell_rsa_0_s0_read),        //               .read
		.avs_s0_write              (mm_interconnect_1_avalon_shell_rsa_0_s0_write),       //               .write
		.avs_s0_readdata           (mm_interconnect_1_avalon_shell_rsa_0_s0_readdata),    //               .readdata
		.avs_s0_writedata          (mm_interconnect_1_avalon_shell_rsa_0_s0_writedata),   //               .writedata
		.avm_design_m0_address     (avalon_shell_rsa_0_m0_address_address),               //     m0_address.address
		.avm_design_m0_read        (avalon_shell_rsa_0_m0_read_read),                     //        m0_read.read
		.avm_design_m0_write       (avalon_shell_rsa_0_m0_write_write),                   //       m0_write.write
		.avm_design_m0_readdata    (avalon_shell_rsa_0_m0_readdata_readdata),             //    m0_readdata.readdata
		.avm_design_m0_writedata   (avalon_shell_rsa_0_m0_writedata_writedata),           //   m0_writedata.writedata
		.avm_design_s0_waitrequest (avalon_shell_rsa_0_s0_waitrequest_waitrequest),       // s0_waitrequest.waitrequest
		.avm_design_s0_address     (avalon_shell_rsa_0_s0_address_address),               //     s0_address.address
		.avm_design_s0_read        (avalon_shell_rsa_0_s0_read_read),                     //        s0_read.read
		.avm_design_s0_write       (avalon_shell_rsa_0_s0_write_write),                   //       s0_write.write
		.avm_design_s0_readdata    (avalon_shell_rsa_0_s0_readdata_readdata),             //    s0_readdata.readdata
		.avm_design_s0_writedata   (avalon_shell_rsa_0_s0_writedata_writedata),           //   s0_writedata.writedata
		.avm_design_m0_waitrequest (avalon_shell_rsa_0_m0_waitrequest_waitrequest)        // m0_waitrequest.waitrequest
	);

	PCIe_rsa_ddr3a ddr3a (
		.pll_ref_clk               (clk_0_clk),                                      //      pll_ref_clk.clk
		.global_reset_n            (reset_0_reset_n),                                //     global_reset.reset_n
		.soft_reset_n              (reset_0_reset_n),                                //       soft_reset.reset_n
		.afi_clk                   (ddr3a_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                               //     afi_half_clk.clk
		.afi_reset_n               (),                                               //        afi_reset.reset_n
		.afi_reset_export_n        (),                                               // afi_reset_export.reset_n
		.mem_a                     (ddr3a_mem_a),                                    //           memory.mem_a
		.mem_ba                    (ddr3a_mem_ba),                                   //                 .mem_ba
		.mem_ck                    (ddr3a_mem_ck),                                   //                 .mem_ck
		.mem_ck_n                  (ddr3a_mem_ck_n),                                 //                 .mem_ck_n
		.mem_cke                   (ddr3a_mem_cke),                                  //                 .mem_cke
		.mem_cs_n                  (ddr3a_mem_cs_n),                                 //                 .mem_cs_n
		.mem_dm                    (ddr3a_mem_dm),                                   //                 .mem_dm
		.mem_ras_n                 (ddr3a_mem_ras_n),                                //                 .mem_ras_n
		.mem_cas_n                 (ddr3a_mem_cas_n),                                //                 .mem_cas_n
		.mem_we_n                  (ddr3a_mem_we_n),                                 //                 .mem_we_n
		.mem_reset_n               (ddr3a_mem_reset_n),                              //                 .mem_reset_n
		.mem_dq                    (ddr3a_mem_dq),                                   //                 .mem_dq
		.mem_dqs                   (ddr3a_mem_dqs),                                  //                 .mem_dqs
		.mem_dqs_n                 (ddr3a_mem_dqs_n),                                //                 .mem_dqs_n
		.mem_odt                   (ddr3a_mem_odt),                                  //                 .mem_odt
		.avl_ready                 (mm_interconnect_2_ddr3a_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_2_ddr3a_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_2_ddr3a_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_2_ddr3a_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_2_ddr3a_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_2_ddr3a_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_2_ddr3a_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_2_ddr3a_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_2_ddr3a_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_2_ddr3a_avl_burstcount),         //                 .burstcount
		.local_init_done           (ddr3a_status_local_init_done),                   //           status.local_init_done
		.local_cal_success         (ddr3a_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail            (ddr3a_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rzqin                 (ddr3a_oct_rzqin),                                //              oct.rzqin
		.pll_mem_clk               (ddr3a_pll_sharing_pll_mem_clk),                  //      pll_sharing.pll_mem_clk
		.pll_write_clk             (ddr3a_pll_sharing_pll_write_clk),                //                 .pll_write_clk
		.pll_locked                (ddr3a_pll_sharing_pll_locked),                   //                 .pll_locked
		.pll_write_clk_pre_phy_clk (ddr3a_pll_sharing_pll_write_clk_pre_phy_clk),    //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (ddr3a_pll_sharing_pll_addr_cmd_clk),             //                 .pll_addr_cmd_clk
		.pll_avl_clk               (ddr3a_pll_sharing_pll_avl_clk),                  //                 .pll_avl_clk
		.pll_config_clk            (ddr3a_pll_sharing_pll_config_clk),               //                 .pll_config_clk
		.pll_hr_clk                (ddr3a_pll_sharing_pll_hr_clk),                   //                 .pll_hr_clk
		.pll_p2c_read_clk          (ddr3a_pll_sharing_pll_p2c_read_clk),             //                 .pll_p2c_read_clk
		.pll_c2p_write_clk         (ddr3a_pll_sharing_pll_c2p_write_clk)             //                 .pll_c2p_write_clk
	);

	PCIe_rsa_dma0 dma0 (
		.clk                (pcie_interface_coreclkout_clk),                        //                clk.clk
		.system_reset_n     (~rst_controller_001_reset_out_reset),                  //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_dma0_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_dma0_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_dma0_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_dma0_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_dma0_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver0_irq),                             //                irq.irq
		.read_address       (dma0_read_master_address),                             //        read_master.address
		.read_chipselect    (dma0_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma0_read_master_read),                                //                   .read_n
		.read_readdata      (dma0_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma0_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma0_read_master_waitrequest),                         //                   .waitrequest
		.read_burstcount    (dma0_read_master_burstcount),                          //                   .burstcount
		.write_address      (dma0_write_master_address),                            //       write_master.address
		.write_chipselect   (dma0_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma0_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma0_write_master_write),                              //                   .write_n
		.write_writedata    (dma0_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma0_write_master_byteenable),                         //                   .byteenable
		.write_burstcount   (dma0_write_master_burstcount)                          //                   .burstcount
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (128),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (10),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) dma0_pp (
		.clk              (pcie_interface_coreclkout_clk),              //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),         // reset.reset
		.s0_waitrequest   (mm_interconnect_3_dma0_pp_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_3_dma0_pp_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_3_dma0_pp_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_3_dma0_pp_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_3_dma0_pp_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_3_dma0_pp_s0_address),       //      .address
		.s0_write         (mm_interconnect_3_dma0_pp_s0_write),         //      .write
		.s0_read          (mm_interconnect_3_dma0_pp_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_3_dma0_pp_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_3_dma0_pp_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (dma0_pp_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (dma0_pp_m0_readdata),                        //      .readdata
		.m0_readdatavalid (dma0_pp_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (dma0_pp_m0_burstcount),                      //      .burstcount
		.m0_writedata     (dma0_pp_m0_writedata),                       //      .writedata
		.m0_address       (dma0_pp_m0_address),                         //      .address
		.m0_write         (dma0_pp_m0_write),                           //      .write
		.m0_read          (dma0_pp_m0_read),                            //      .read
		.m0_byteenable    (dma0_pp_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (dma0_pp_m0_debugaccess)                      //      .debugaccess
	);

	PCIe_rsa_mm_interconnect_0 mm_interconnect_0 (
		.PCIE_interface_coreclkout_clk          (pcie_interface_coreclkout_clk),                        //        PCIE_interface_coreclkout.clk
		.dma0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                   // dma0_reset_reset_bridge_in_reset.reset
		.PCIE_interface_Rxm_BAR0_address        (pcie_interface_rxm_bar0_address),                      //          PCIE_interface_Rxm_BAR0.address
		.PCIE_interface_Rxm_BAR0_waitrequest    (pcie_interface_rxm_bar0_waitrequest),                  //                                 .waitrequest
		.PCIE_interface_Rxm_BAR0_burstcount     (pcie_interface_rxm_bar0_burstcount),                   //                                 .burstcount
		.PCIE_interface_Rxm_BAR0_byteenable     (pcie_interface_rxm_bar0_byteenable),                   //                                 .byteenable
		.PCIE_interface_Rxm_BAR0_read           (pcie_interface_rxm_bar0_read),                         //                                 .read
		.PCIE_interface_Rxm_BAR0_readdata       (pcie_interface_rxm_bar0_readdata),                     //                                 .readdata
		.PCIE_interface_Rxm_BAR0_readdatavalid  (pcie_interface_rxm_bar0_readdatavalid),                //                                 .readdatavalid
		.PCIE_interface_Rxm_BAR0_write          (pcie_interface_rxm_bar0_write),                        //                                 .write
		.PCIE_interface_Rxm_BAR0_writedata      (pcie_interface_rxm_bar0_writedata),                    //                                 .writedata
		.dma0_control_port_slave_address        (mm_interconnect_0_dma0_control_port_slave_address),    //          dma0_control_port_slave.address
		.dma0_control_port_slave_write          (mm_interconnect_0_dma0_control_port_slave_write),      //                                 .write
		.dma0_control_port_slave_readdata       (mm_interconnect_0_dma0_control_port_slave_readdata),   //                                 .readdata
		.dma0_control_port_slave_writedata      (mm_interconnect_0_dma0_control_port_slave_writedata),  //                                 .writedata
		.dma0_control_port_slave_chipselect     (mm_interconnect_0_dma0_control_port_slave_chipselect), //                                 .chipselect
		.PCIE_interface_Cra_address             (mm_interconnect_0_pcie_interface_cra_address),         //               PCIE_interface_Cra.address
		.PCIE_interface_Cra_write               (mm_interconnect_0_pcie_interface_cra_write),           //                                 .write
		.PCIE_interface_Cra_read                (mm_interconnect_0_pcie_interface_cra_read),            //                                 .read
		.PCIE_interface_Cra_readdata            (mm_interconnect_0_pcie_interface_cra_readdata),        //                                 .readdata
		.PCIE_interface_Cra_writedata           (mm_interconnect_0_pcie_interface_cra_writedata),       //                                 .writedata
		.PCIE_interface_Cra_byteenable          (mm_interconnect_0_pcie_interface_cra_byteenable),      //                                 .byteenable
		.PCIE_interface_Cra_waitrequest         (mm_interconnect_0_pcie_interface_cra_waitrequest),     //                                 .waitrequest
		.PCIE_interface_Cra_chipselect          (mm_interconnect_0_pcie_interface_cra_chipselect)       //                                 .chipselect
	);

	PCIe_rsa_mm_interconnect_1 mm_interconnect_1 (
		.clk_clk_clk                                                          (clk_0_clk),                                           //                                                        clk_clk.clk
		.PCIE_interface_coreclkout_clk                                        (pcie_interface_coreclkout_clk),                       //                                      PCIE_interface_coreclkout.clk
		.avalon_shell_rsa_0_reset_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                      //                 avalon_shell_rsa_0_reset_reset_bridge_in_reset.reset
		.PCIE_interface_Rxm_BAR2_translator_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                  // PCIE_interface_Rxm_BAR2_translator_reset_reset_bridge_in_reset.reset
		.PCIE_interface_Rxm_BAR2_address                                      (pcie_interface_rxm_bar2_address),                     //                                        PCIE_interface_Rxm_BAR2.address
		.PCIE_interface_Rxm_BAR2_waitrequest                                  (pcie_interface_rxm_bar2_waitrequest),                 //                                                               .waitrequest
		.PCIE_interface_Rxm_BAR2_burstcount                                   (pcie_interface_rxm_bar2_burstcount),                  //                                                               .burstcount
		.PCIE_interface_Rxm_BAR2_byteenable                                   (pcie_interface_rxm_bar2_byteenable),                  //                                                               .byteenable
		.PCIE_interface_Rxm_BAR2_read                                         (pcie_interface_rxm_bar2_read),                        //                                                               .read
		.PCIE_interface_Rxm_BAR2_readdata                                     (pcie_interface_rxm_bar2_readdata),                    //                                                               .readdata
		.PCIE_interface_Rxm_BAR2_readdatavalid                                (pcie_interface_rxm_bar2_readdatavalid),               //                                                               .readdatavalid
		.PCIE_interface_Rxm_BAR2_write                                        (pcie_interface_rxm_bar2_write),                       //                                                               .write
		.PCIE_interface_Rxm_BAR2_writedata                                    (pcie_interface_rxm_bar2_writedata),                   //                                                               .writedata
		.avalon_shell_rsa_0_s0_address                                        (mm_interconnect_1_avalon_shell_rsa_0_s0_address),     //                                          avalon_shell_rsa_0_s0.address
		.avalon_shell_rsa_0_s0_write                                          (mm_interconnect_1_avalon_shell_rsa_0_s0_write),       //                                                               .write
		.avalon_shell_rsa_0_s0_read                                           (mm_interconnect_1_avalon_shell_rsa_0_s0_read),        //                                                               .read
		.avalon_shell_rsa_0_s0_readdata                                       (mm_interconnect_1_avalon_shell_rsa_0_s0_readdata),    //                                                               .readdata
		.avalon_shell_rsa_0_s0_writedata                                      (mm_interconnect_1_avalon_shell_rsa_0_s0_writedata),   //                                                               .writedata
		.avalon_shell_rsa_0_s0_waitrequest                                    (mm_interconnect_1_avalon_shell_rsa_0_s0_waitrequest)  //                                                               .waitrequest
	);

	PCIe_rsa_mm_interconnect_2 mm_interconnect_2 (
		.clk_clk_clk                                            (clk_0_clk),                                          //                                          clk_clk.clk
		.ddr3a_afi_clk_clk                                      (ddr3a_afi_clk_clk),                                  //                                    ddr3a_afi_clk.clk
		.PCIE_interface_coreclkout_clk                          (pcie_interface_coreclkout_clk),                      //                        PCIE_interface_coreclkout.clk
		.avalon_shell_rsa_0_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                     //   avalon_shell_rsa_0_reset_reset_bridge_in_reset.reset
		.ddr3a_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                 // ddr3a_avl_translator_reset_reset_bridge_in_reset.reset
		.ddr3a_soft_reset_reset_bridge_in_reset_reset           (rst_controller_002_reset_out_reset),                 //           ddr3a_soft_reset_reset_bridge_in_reset.reset
		.dma0_pp_reset_reset_bridge_in_reset_reset              (rst_controller_001_reset_out_reset),                 //              dma0_pp_reset_reset_bridge_in_reset.reset
		.avalon_shell_rsa_0_m0_address                          (avalon_shell_rsa_0_m0_address),                      //                            avalon_shell_rsa_0_m0.address
		.avalon_shell_rsa_0_m0_waitrequest                      (avalon_shell_rsa_0_m0_waitrequest),                  //                                                 .waitrequest
		.avalon_shell_rsa_0_m0_read                             (avalon_shell_rsa_0_m0_read),                         //                                                 .read
		.avalon_shell_rsa_0_m0_readdata                         (avalon_shell_rsa_0_m0_readdata),                     //                                                 .readdata
		.avalon_shell_rsa_0_m0_write                            (avalon_shell_rsa_0_m0_write),                        //                                                 .write
		.avalon_shell_rsa_0_m0_writedata                        (avalon_shell_rsa_0_m0_writedata),                    //                                                 .writedata
		.dma0_pp_m0_address                                     (dma0_pp_m0_address),                                 //                                       dma0_pp_m0.address
		.dma0_pp_m0_waitrequest                                 (dma0_pp_m0_waitrequest),                             //                                                 .waitrequest
		.dma0_pp_m0_burstcount                                  (dma0_pp_m0_burstcount),                              //                                                 .burstcount
		.dma0_pp_m0_byteenable                                  (dma0_pp_m0_byteenable),                              //                                                 .byteenable
		.dma0_pp_m0_read                                        (dma0_pp_m0_read),                                    //                                                 .read
		.dma0_pp_m0_readdata                                    (dma0_pp_m0_readdata),                                //                                                 .readdata
		.dma0_pp_m0_readdatavalid                               (dma0_pp_m0_readdatavalid),                           //                                                 .readdatavalid
		.dma0_pp_m0_write                                       (dma0_pp_m0_write),                                   //                                                 .write
		.dma0_pp_m0_writedata                                   (dma0_pp_m0_writedata),                               //                                                 .writedata
		.dma0_pp_m0_debugaccess                                 (dma0_pp_m0_debugaccess),                             //                                                 .debugaccess
		.ddr3a_avl_address                                      (mm_interconnect_2_ddr3a_avl_address),                //                                        ddr3a_avl.address
		.ddr3a_avl_write                                        (mm_interconnect_2_ddr3a_avl_write),                  //                                                 .write
		.ddr3a_avl_read                                         (mm_interconnect_2_ddr3a_avl_read),                   //                                                 .read
		.ddr3a_avl_readdata                                     (mm_interconnect_2_ddr3a_avl_readdata),               //                                                 .readdata
		.ddr3a_avl_writedata                                    (mm_interconnect_2_ddr3a_avl_writedata),              //                                                 .writedata
		.ddr3a_avl_beginbursttransfer                           (mm_interconnect_2_ddr3a_avl_beginbursttransfer),     //                                                 .beginbursttransfer
		.ddr3a_avl_burstcount                                   (mm_interconnect_2_ddr3a_avl_burstcount),             //                                                 .burstcount
		.ddr3a_avl_byteenable                                   (mm_interconnect_2_ddr3a_avl_byteenable),             //                                                 .byteenable
		.ddr3a_avl_readdatavalid                                (mm_interconnect_2_ddr3a_avl_readdatavalid),          //                                                 .readdatavalid
		.ddr3a_avl_waitrequest                                  (~mm_interconnect_2_ddr3a_avl_waitrequest),           //                                                 .waitrequest
		.PCIE_interface_Txs_address                             (mm_interconnect_2_pcie_interface_txs_address),       //                               PCIE_interface_Txs.address
		.PCIE_interface_Txs_write                               (mm_interconnect_2_pcie_interface_txs_write),         //                                                 .write
		.PCIE_interface_Txs_read                                (mm_interconnect_2_pcie_interface_txs_read),          //                                                 .read
		.PCIE_interface_Txs_readdata                            (mm_interconnect_2_pcie_interface_txs_readdata),      //                                                 .readdata
		.PCIE_interface_Txs_writedata                           (mm_interconnect_2_pcie_interface_txs_writedata),     //                                                 .writedata
		.PCIE_interface_Txs_burstcount                          (mm_interconnect_2_pcie_interface_txs_burstcount),    //                                                 .burstcount
		.PCIE_interface_Txs_byteenable                          (mm_interconnect_2_pcie_interface_txs_byteenable),    //                                                 .byteenable
		.PCIE_interface_Txs_readdatavalid                       (mm_interconnect_2_pcie_interface_txs_readdatavalid), //                                                 .readdatavalid
		.PCIE_interface_Txs_waitrequest                         (mm_interconnect_2_pcie_interface_txs_waitrequest),   //                                                 .waitrequest
		.PCIE_interface_Txs_chipselect                          (mm_interconnect_2_pcie_interface_txs_chipselect)     //                                                 .chipselect
	);

	PCIe_rsa_mm_interconnect_3 mm_interconnect_3 (
		.PCIE_interface_coreclkout_clk          (pcie_interface_coreclkout_clk),              //        PCIE_interface_coreclkout.clk
		.dma0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),         // dma0_reset_reset_bridge_in_reset.reset
		.dma0_read_master_address               (dma0_read_master_address),                   //                 dma0_read_master.address
		.dma0_read_master_waitrequest           (dma0_read_master_waitrequest),               //                                 .waitrequest
		.dma0_read_master_burstcount            (dma0_read_master_burstcount),                //                                 .burstcount
		.dma0_read_master_chipselect            (dma0_read_master_chipselect),                //                                 .chipselect
		.dma0_read_master_read                  (~dma0_read_master_read),                     //                                 .read
		.dma0_read_master_readdata              (dma0_read_master_readdata),                  //                                 .readdata
		.dma0_read_master_readdatavalid         (dma0_read_master_readdatavalid),             //                                 .readdatavalid
		.dma0_write_master_address              (dma0_write_master_address),                  //                dma0_write_master.address
		.dma0_write_master_waitrequest          (dma0_write_master_waitrequest),              //                                 .waitrequest
		.dma0_write_master_burstcount           (dma0_write_master_burstcount),               //                                 .burstcount
		.dma0_write_master_byteenable           (dma0_write_master_byteenable),               //                                 .byteenable
		.dma0_write_master_chipselect           (dma0_write_master_chipselect),               //                                 .chipselect
		.dma0_write_master_write                (~dma0_write_master_write),                   //                                 .write
		.dma0_write_master_writedata            (dma0_write_master_writedata),                //                                 .writedata
		.dma0_pp_s0_address                     (mm_interconnect_3_dma0_pp_s0_address),       //                       dma0_pp_s0.address
		.dma0_pp_s0_write                       (mm_interconnect_3_dma0_pp_s0_write),         //                                 .write
		.dma0_pp_s0_read                        (mm_interconnect_3_dma0_pp_s0_read),          //                                 .read
		.dma0_pp_s0_readdata                    (mm_interconnect_3_dma0_pp_s0_readdata),      //                                 .readdata
		.dma0_pp_s0_writedata                   (mm_interconnect_3_dma0_pp_s0_writedata),     //                                 .writedata
		.dma0_pp_s0_burstcount                  (mm_interconnect_3_dma0_pp_s0_burstcount),    //                                 .burstcount
		.dma0_pp_s0_byteenable                  (mm_interconnect_3_dma0_pp_s0_byteenable),    //                                 .byteenable
		.dma0_pp_s0_readdatavalid               (mm_interconnect_3_dma0_pp_s0_readdatavalid), //                                 .readdatavalid
		.dma0_pp_s0_waitrequest                 (mm_interconnect_3_dma0_pp_s0_waitrequest),   //                                 .waitrequest
		.dma0_pp_s0_debugaccess                 (mm_interconnect_3_dma0_pp_s0_debugaccess)    //                                 .debugaccess
	);

	PCIe_rsa_irq_mapper irq_mapper (
		.clk           (pcie_interface_coreclkout_clk),      //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (pcie_interface_rxmirq_irq)           //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_0_reset_n),               // reset_in0.reset
		.clk            (clk_0_clk),                      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~pcie_interface_nreset_status_reset), // reset_in0.reset
		.clk            (pcie_interface_coreclkout_clk),       //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_in1      (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_0_reset_n),                   // reset_in0.reset
		.clk            (ddr3a_afi_clk_clk),                  //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
